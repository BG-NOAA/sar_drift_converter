netcdf SAR_drift_data {
dimensions:
	time = UNLIMITED ; // (0 currently)
	y = 361 ;
	x = 361 ;
variables:
	float Speed_kmdy(time, y, x) ;
		Speed_kmdy:long_name = "Speed in km/day" ;
		Speed_kmdy:standard_name = "sea_ice_speed" ;
		Speed_kmdy:ioos_category = "SAR daily sea-ice drift" ;
		Speed_kmdy:units = "km/day" ;
		Speed_kmdy:grid_mapping = "spatial_ref" ;
	float dx(time, y, x) ;
		dx:_FillValue = NaNf ;
		dx:long_name = "Zonal Velocity" ;
		dx:standard_name = "movement_in_x_direction" ;
		dx:ioos_category = "SAR daily sea-ice drift" ;
		dx:units = "m/day" ;
		dx:grid_mapping = "spatial_ref" ;
	float dy(time, y, x) ;
		dy:_FillValue = NaNf ;
		dy:long_name = "Meridional Velocity" ;
		dy:standard_name = "movement_in_y_direction" ;
		dy:ioos_category = "SAR daily sea-ice drift" ;
		dy:units = "m/day" ;
		dy:grid_mapping = "spatial_ref" ;
	float Bear_deg(time, y, x) ;
		Bear_deg:long_name = "Bearing" ;
		Bear_deg:standard_name = "direction_true_north" ;
		Bear_deg:ioos_category = "SAR daily sea-ice drift" ;
		Bear_deg:units = "degrees" ;
		Bear_deg:grid_mapping = "spatial_ref" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Centered Time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double x(x) ;
		x:standard_name = "projection_x_coordinate" ;
		x:long_name = "x coordinate of projection" ;
		x:units = "m" ;
		x:axis = "X" ;
	double y(y) ;
		y:standard_name = "projection_y_coordinate" ;
		y:long_name = "y coordinate of projection" ;
		y:units = "m" ;
		y:axis = "Y" ;
	int spatial_ref ;
		spatial_ref:grid_mapping_name = "polar_stereographic" ;
		spatial_ref:straight_vertical_longitude_from_pole = -45. ;
		spatial_ref:latitude_of_projection_origin = 90. ;
		spatial_ref:standard_parallel = 70. ;
		spatial_ref:false_easting = 0. ;
		spatial_ref:false_northing = 0. ;
		spatial_ref:semi_major_axis = 6378137. ;
		spatial_ref:inverse_flattening = 298.2794111 ;
		spatial_ref:spatial_ref = "EPSG:3413" ;
		spatial_ref:crs = "PROJCS[\"WGS 84 / NSIDC Sea Ice Polar Stereographic North\",GEOGCS[\"WGS 84\",DATUM[\"WGS_1984\",SPHEROID[\"WGS 84\",6378137,298.257223563]],PRIMEM[\"Greenwich\",0],UNIT[\"degree\",0.0174532925199433]],PROJECTION[\"Polar_Stereographic\"],PARAMETER[\"latitude_of_origin\",70],PARAMETER[\"central_meridian\",-45],PARAMETER[\"scale_factor\",1],PARAMETER[\"false_easting\",0],PARAMETER[\"false_northing\",0],UNIT[\"metre\",1,AUTHORITY[\"EPSG\",\"9001\"]]]" ;

// global attributes:
		:Conventions = "CF-1.8, ACDD-1.3" ;
		:title = "SAR drift data converted from raw text form to NetCDF" ;
		:summary = "NetCDF version of the SAR Daily Drift dataset. This dataset includes the starting and ending coordinates (latitude and longitude), start and end observation dates, total distance traveled, and drift bearing over the observation period." ;
		:acknowledgement = "Produced by NOAA using IABP data." ;
		:creator_name = "Brendon Gory" ;
		:creator_email = "brendon.gory@noaa.gov" ;
		:creator_institution = "CIRA/NOAA" ;
		:creator_type = "Institution" ;
		:creator_url = "https://noaa.gov/" ;
		:publisher_name = "NOAA CoastWatch" ;
		:publisher_email = "coastwatch@noaa.gov" ;
		:publisher_institution = "NOAA CoastWatch" ;
		:publisher_type = "Institutional" ;
		:publisher_url = "https://coastwatch.noaa.gov/" ;
		:contributor_name = "NOAA PolarWatch, Southwest Fisheries Science Center, NESDIS STAR, U.S. National Ice Center" ;
		:contributor_role = "Producer, Publisher, Advisor, Originator" ;
		:processing_level = "NOAA Level 4" ;
		:product_version = "Version 1" ;
		:project = "NOAA Polarwatch" ;
		:source = "SAR Daily Drift dataset" ;
		:instrument = "See website for details" ;
		:platform = "Earth Observation Satellites, In Situ Land-based Platforms, Ground Stations, Models/Analyses" ;
		:platform_vocabulary = "NASA Global Change Master Directory (GCMD) Keywords, Version 9.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (Version 72, 10 March 2020)" ;
		:keywords = "Earth Science > Cryosphere > Sea Ice > Ice Extent, Earth Science > Cryosphere > Snow/Ice > Snow Cover, GEOGRAPHIC REGION > ARCTIC, GEOGRAPHIC REGION > NORTHERN HEMISPHERE, GEOGRAPHIC REGION > POLAR" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Keywords, Version 9.0" ;
		:license = "U.S. Government Work (public domain)" ;
		:history = "2025-04-02: First version of convert SAR daily drift to NetCDF" ;
		:references = "https://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
		:metadata_link = "https://coastwatch.noaa.gov/cwn/products/sar-composite-arctic-imagery-normalized-radar-cross-section.html" ;
		:sourceUrl = "https://www.star.nesdis.noaa.gov/socd/mecb/sar/AKDEMO_products/COMPOSITE_TIFF/DRIFT_SHAPEFILES/" ;
		:naming_authority = "gov.noaa.polarwatch" ;
		:ncei_template_version = "NCEI_NetCDF_Grid_Template_v2.0" ;
		:date_created = "FILL_DATE_CREATED" ;
		:time_coverage_start = "FILL_MIN_TIME" ;
		:time_coverage_end = "FILL_MAX_TIME" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_resolution = "P1D" ;
}